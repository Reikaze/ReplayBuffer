`include "crc.v"

module crc_tb;

reg clk_t;
reg rst_t;
reg we_t;
reg [27:0] tlp_in_t;

wire [15:0] crc_out_t;






endmodule
